
.MODEL PX1 PNP (RB = 163.5 IRB = 0 RBM = 12.27 RC = 25 RE = 1.5
+ IS = 147E-18 EG = 1.206 XTI = 1.7 XTB = 1.866 BF = 110.0
+ IKF = 4.718E-3 NF = 1 VAF = 51.8 ISE = 50.2E-16 NE = 1.65
+ BR = 0.4745 IKR = 12.96E-3 NR = 1 VAR = 9.96 ISC = 0 NC = 2
+ TF = 0.610E-9 TR = 0.610E-8 CJE = 0.36E-12 VJE = 0.5
+ MJE = 0.28 CJC = 0.328E-12 VJC = 0.8 MJC = 0.4 XCJC = 0.074
+ CJS = 1.39E-12 VJS = 0.55 MJS = 0.35 FC = 0.5)

.MODEL NX1 NPN (RB = 262.5 IRB = 0 RBM = 12.5 RC = 25 RE = 0.5
+ IS = 242E-18 EG = 1.206 XTI = 2 XTB = 1.538 BF = 137.5
+ IKF = 13.94E-3 NF = 1.0 VAF = 159.4 ISE = 72E-16 NE = 1.713
+ BR = 0.7258 IKR = 4.396E-3 NR = 1.0 VAR = 10.73 ISC = 0 NC = 2
+ TF = 0.425E-9 TR = 0.425E-8 CJE = 0.428E-12 VJE = 0.5
+ MJE = 0.28 CJC = 1.97E-13 VJC = 0.5 MJC = 0.3 XCJC = 0.065
+ CJS = 1.17E-12 VJS = 0.64 MJS = 0.4 FC = 0.5)

Q1 8 8 0 NX1
Q2 7 7 8 NX1
Q3 1 7 6 NX1
Q4 5 6 0 NX1
Q5 2 3 0 NX1
Q6 3 3 0 NX1

Q7 2 2 1 PX1
Q8 8 2 1 PX1
Q9 5 5 1 PX1
Q10 4 5 1 PX1
Q11 10 5 1 PX1

If1 1 7 50uA
If2 8 0 50uA
If3 6 0 50uA
Iu 4 3 ac 20uA

Vlp 10 11 0V
Vhp 4 11 0V

RL 11 0 1

C1 6 0 300pF

VCC 1 0 3V


*.DC Iu 10uA 40uA 0.01uA
.AC dec 100 1 10meg