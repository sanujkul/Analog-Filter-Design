*Following is circuit implementation of LP, HP, BP filters from
*a two CFOAs
* based on Lab Experiment 8 in course ECD07
* by Prof. Raj Senani

.include /Users/sanujkul/Documents/LTspice/libraries/ad844.cir
*i. CFOAs:
*Xn Y X +V -V W Z MODELNAME
X1 3 2 7 4 6 5 AD844
X2 6 8 7 4 10 9 AD844

*ii. Passive Componets
R1 1 8 707
R2 9 0 707
R3 3 10 1.41k
C1 5 0 1n
C2 9 11 1n

*iii. Power supplies:
VccPositive 7 0 DC 12V
VccNegative 4 0 DC -12V

*iv. Voltage inputs:
*LP: V2=V3=0, BP: V1=V3=0, HP:V2=V1=0
*AP: V1=V2=V3, R1=R2, BR: V2=0
V1 2 0 AC 1mV
V2 1 0 AC 0mv
V3 11 0 AC 0mV

***** OUTPUT CODES **********
*AC ANALYSIS
.AC DEC 50 10K 20MEG
***************************************
*Nwxt two lines for TRANSIENT ANALYSIS
*VT 2 0 PULSE(0 1.8 0 1n 1n 10n 22n)
*.tran 0 100n
***************************************
*DC ANALYSIS
*VT 2 0 DC 1V
*.dc Vt 0 1.8 0.1
***************************************

