*Following is circuit implementation of LP, HP, BP filters from
*a two CFOAs
* based on Lab Experiment 8 in course ECD07
* by Prof. Raj Senani

.include /Users/sanujkul/Documents/LTspice/Workspace/Analog-Filter-Design/Exp09-Tunable-BP-CCII/CCII-subckt/CCII.cir
*CCIIs:
*.SUBCKT CCIIplus Y X Z Vdd Vss Ib
XCCii1 1 2 4 100 101 3 CCIIplus
XCCii2 5 4 7 100 101 6 CCIIplus
XCCii3 7 8 4 100 101 9 CCIIplus

*Capacitors:
C1 7 0 50p
C2 4 0 50p

*VOLTAGE SOURCES:
Vdd 100 0 DC 12V
Vss 101 0 DC -12V

Vin 1 0 AC 1mV
Vx1 2 0 DC 0V
Vy2 5 0 DC 0V
Vx3 8 0 DC 0V

*CURRENT SOURCES:
Ib1 0 3 DC 0.5mA
Ib2 0 6 DC 0.5mA
Ib3 0 9 DC {values3}
.param values3 = 1
.step param values3 list 0.1uA 10uA 100uA 1mA


***** OUTPUT CODES **********
*AC ANALYSIS
.AC DEC 50 1K 10G
***************************************
*Nwxt two lines for TRANSIENT ANALYSIS
*VT 2 0 PULSE(0 1.8 0 1n 1n 10n 22n)
*.tran 0 100n
***************************************
*DC ANALYSIS
*VT 2 0 DC 1V
*.dc Vt 0 1.8 0.1
***************************************

